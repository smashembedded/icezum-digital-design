// Baud generator
`include "../baudgen/baudgen_tx.v"