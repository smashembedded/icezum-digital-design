//-------------------------------------------------------------------
//-- or4.v
//-- Module
//-------------------------------------------------------------------
//-- Daniel Rodrigo
//-- GPL license
//-------------------------------------------------------------------
//-- OR Logic Gate 4:1
//-------------------------------------------------------------------

module or4 (x0, x1, x2, x3, z0);

// inputs and output
input x0, x1, x2, x3;
output z0;

// define signals
wire x0, x1, x2, x3;
wire z0;

// continuous assign
assign z0 = x0 | x1 | x2 | x3;

endmodule