// Baud generator
`include "../baudgen/baudgen_rx.v"