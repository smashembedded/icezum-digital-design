//-------------------------------------------------------------------
//-- and2.v
//-- Testbench
//-------------------------------------------------------------------
//-- Daniel Rodrigo
//-- GPL license
//-------------------------------------------------------------------

module and2 (SW1, SW2, LED0);

input SW1, SW2;
output LED0;

wire SW1, SW2;
wire LED0;

assign LED0 = SW1 & SW2;

endmodule